`timescale 1ns/1ps

module UART_Rx #(parameter UART_CLK_FREQ = 150_000_000,   // UART Input Clock Frequency
                          BAUD_RATE = 3_000_000,        // Desired Baud Rate
                          OVERSAMPLING = 16            // Oversampling factor (default is 16×)
)(
    //input wire CLK,         // System clock input (e.g., 150 MHz)
    input wire BCLK,
    input wire RST,         // Active-high synchronous reset
    input wire RX,          // UART receive signal

    //output reg [7:0] RDATA, // Received data
    output reg [7:0] DOUT,
    output reg DONERX       // Receive complete signal
);

    // Internal signals
   // wire BCLK;              // Baud clock generated by baud_gen module
    reg [7:0] RDATA;

    // Instantiate the baud rate generator
   /* baud_gen #(
        .UART_CLK_FREQ(UART_CLK_FREQ),
        .BAUD_RATE(BAUD_RATE),
        .OVERSAMPLING(OVERSAMPLING)
    ) baud_gen_inst (
        .CLK(CLK),          // System clock input
        .RST(RST),          // Active-high reset
        .BCLK(BCLK)         // Generated baud clock output
    ); */

    // State encoding
    localparam IDLE = 2'b00, START = 2'b01, END = 2'b10;

    // Registers
    reg [1:0]pr_state;           // Present state
    reg [3:0] counts;       // Bit counter for receiving data (0 to 7)

    // State machine
    always @(posedge BCLK or posedge RST) begin
        if (RST) begin
            pr_state <= IDLE;
            DOUT <= 8'b0;
            RDATA <= 8'b0;
            DONERX <= 1'b0;
            counts <= 4'd0;
        end else begin
            case (pr_state)
                IDLE: begin
                    DONERX <= 1'b0;   // Clear receive complete flag
                    RDATA <= 8'b0;    // Clear data register
                    if (RX == 1'b0) begin
                        pr_state <= START; // Start bit detected
                    end else begin
                        pr_state <= IDLE;
                    end
                end

                START: begin
                    if (counts < 8) begin
                        RDATA <= {RDATA[6:0], RX}; // Shift in received bit
                        counts <= counts + 1;
                        pr_state <= START;
                    end else begin
                        DONERX <= 1'b1; // Set receive complete flag
                        counts <= 4'd0; // Reset bit counter
                        DOUT <= RDATA;
                        pr_state <= END;
                    end
                end
                
                END: begin
                    if(DONERX == 1)begin
                       // DOUT <= RDATA;
                        DONERX <= 0;
                    end
                    pr_state <= IDLE;
                end

                default: pr_state <= IDLE; // Default state
            endcase
        end
    end

endmodule