`timescale 1ns/1ps

module UART_Tx #(parameter UART_CLK_FREQ = 150_000_000,   // UART Input Clock Frequency
                          BAUD_RATE = 3_000_000,        // Desired Baud Rate
                          OVERSAMPLING = 16            // Oversampling factor (default is 16×)
)(
    //input wire CLK,         // System clock input (e.g., 150 MHz)
    input wire BCLK,
    input wire RST,         // Active-high synchronous reset
    input wire NEWD,        // New data signal
    input wire [7:0] TDATA, // Data to transmit

    output reg TX,          // UART transmit signal
    output reg DONETX       // Transmit done signal
);

    // Internal signals
    //wire BCLK;              // Baud clock generated by baud_gen module

    // Instantiate the baud rate generator
    /*baud_gen #(
        .UART_CLK_FREQ(UART_CLK_FREQ),
        .BAUD_RATE(BAUD_RATE),
        .OVERSAMPLING(OVERSAMPLING)
    ) baud_gen_inst (
        .CLK(CLK),          // System clock input
        .RST(RST),          // Active-high reset
        .BCLK(BCLK)         // Generated baud clock output
    ); */

    // State encoding
    localparam [1:0] IDLE = 2'b00, START = 2'b01, TRANS = 2'b10, DONE = 2'b11;

    // Registers
    reg [1:0] pr_state;      // Present state
    reg [3:0] counts;        // Bit counter for transmission (0 to 7)

    // State machine
    always @(posedge BCLK or posedge RST) begin
        if (RST) begin
            pr_state <= IDLE;
            TX <= 1'b1;           // UART line idle (high state)
            DONETX <= 1'b0;
            counts <= 4'd0;
        end else begin
            case (pr_state)
                IDLE: begin
                    TX <= 1'b1;   // UART line idle (high state)
                    DONETX <= 1'b0;
                    if (NEWD) begin
                        pr_state <= START;
                    end else begin
                        pr_state <= IDLE;
                    end
                end

                START: begin
                    TX <= 1'b0;   // Start bit (low state)
                    counts <= 4'b0; // Reset bit counter
                    pr_state <= TRANS;
                    
                end

                TRANS: begin
                    if (counts < 8) begin
                        TX <= TDATA[counts]; // Transmit data bits (LSB first)
                        counts <= counts + 1;
                        pr_state <= TRANS;
                    end else begin
                        TX <= 1'b1; // Stop bit (high state)
                        if(counts == 8)begin
                        DONETX <= 1'b1;
                        end
                        pr_state <= DONE;
                    end
                end

                DONE: begin
               // if(counts == 8)
                    //DONETX <= 1'b1; // Indicate transmission complete
                    pr_state <= IDLE;
                end

                default: pr_state <= IDLE; // Default state
            endcase
        end
    end

endmodule